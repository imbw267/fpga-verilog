//Experiment X
//Author: Brian X. Wu
//Chapter X
//Page X
//Copyright 2017

// Simulation time scale of 1ns
// timestep of 10 ps

`timescale 1 ns/ 10ps

module template_tb();

    // test signal declaration
    localparam T=20;
    wire clk, reset;
    wire data;
    wire dout;

    // instantiate devices under test
    
    // instantiate test vector generator
    // clock is generated here
    

    // instantiate test monitor
    


endmodule