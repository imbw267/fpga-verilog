//Listing 1.3
//Author: Pong P. Chu
//Chapter 1
//Page 8
//Copyright 2008

module eq2_sop
    (
    input wire[1:0] a,b,
    output wire aeqb
    );
    
    // internal signal declaration
    wire p0, p1, p2, p3
    
    // sum of product terms
    assign aeqb = p0 | p1 | p2 | p3;
    
    // product terms
    assign p0 = (~a[1] & ~b[1]) & (~a[0] & ~b[0]);
    assign p1 = (~a[1] & ~b[1]) & (a[0] & b[0]);
    assign p2 = (a[1] & b[1]) & (~a[0] & ~b[0]);
    assign p3 = (a[1] & b[1]) & (a[0] & b[0]);
    
endmodule;  // eq2_sop
     