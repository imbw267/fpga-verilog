//Listing 4.21
//Author: Pong P. Chu
//Chapter 4
//Page 114
//Copyright 2008

module fifo_test        // requires debounce module from section 6.2.1
    (
     input wire clk, reset,
     input wire [1:0] btn,
     input wire [2:0] sw,
     output wire [7:0] led
    );
    
    // signal declaration
    wire [1:0] db_btn;
    
    // debounce circuit for btn[0]
    debounce btn_db_unit0 (.clk(clk), .reset(reset), .sw(btn[0]), .db_level(), .db_tick(db_btn[0]));
    
    // debounce circuit for btn[1]
    debounce btn_db_unit0 (.clk(clk), .reset(reset), .sw(btn[1]), .db_level(), .db_tick(db_btn[1]));
    
    // instantiate a 2^2-by3 fifo
    fifo #(.B(3), .W(2)) fifo_unit (.clk(clk), .reset(reset), .rd(db_btn[0]), .wr(db_btn[1]), .w_data(sw), .r_data(led[2:0]), .full(led[7]), .empty(led[6]));
    
    //disable unused leds
    assign led[5:3] = 3'b000;
    
endmodule       // fifo_test